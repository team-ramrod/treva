--
--  Copyright 2011 Martin Schoeberl <masca@imm.dtu.dk>,
--                 Technical University of Denmark, DTU Informatics. 
--  All rights reserved.
--
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions are met:
-- 
--    1. Redistributions of source code must retain the above copyright notice,
--       this list of conditions and the following disclaimer.
-- 
--    2. Redistributions in binary form must reproduce the above copyright
--       notice, this list of conditions and the following disclaimer in the
--       documentation and/or other materials provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDER ``AS IS'' AND ANY EXPRESS
-- OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES
-- OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED. IN
-- NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE FOR ANY
-- DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
-- LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND
-- ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
-- (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF
-- THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation are
-- those of the authors and should not be interpreted as representing official
-- policies, either expressed or implied, of the copyright holder.
-- 

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.leros_types.all;

-- Some fmax number with Cyclone EP1C12C6
--
--	Memory is with rdaddr in clock process, rddata combinational
--		which is the 'normal' memory configuration, but Quartus
--		adds path through logic for read during write
--	fully registered on-chip memory 256 MHz
--	only input registers, output goes to a LC register (with reset): 165 MHz
--	plus a 16-bit adder: 147 MHz
--	more in ALU + opd mux: 135 MHz
--
--	Memory with rddata in clock process, rdaddr combinational
--		what does this model in read during write? Probably the
--		old value.
--	only input registers, output goes to a LC register (with reset): 256 MHz
--	plus a 16-bit adder: 166 MHz
--	more in ALU (add/sub) and opd mux between imm and DM output: 148 MHz


entity leros_ex is
	port  (
		clk : in std_logic;
		reset : in std_logic;
		din : in fedec_out_type;
		ioin : in io_in_type;
		dout : out ex_out_type
	);
end leros_ex;

architecture rtl of leros_ex is

	-- the accu
	signal accu, opd  : stream_unsigned;
	signal log, arith, a_mux : stream_unsigned;
	
	-- the data ram
	constant nwords : integer := 2 ** DM_BITS;
	type ram_type is array(0 to nwords-1) of std_logic_vector(15 downto 0);
	type ram_array_type is array(0 to stream-1) of ram_type;

	-- 0 initialization is for simulation only
	-- Xilinx and Altera FPGA initialize memory blocks to 0
	signal dm : ram_array_type := (others => (others => (others => '0')));
	
	signal wrdata, rddata : stream_std;
	signal wraddr, rdaddr : std_logic_vector(DM_BITS-1 downto 0);
	
	signal wraddr_dly : std_logic_vector(DM_BITS-1 downto 0);
	signal pc_dly : std_logic_vector(IM_BITS-1 downto 0);
	

begin

	dout.accu <= std_logic_vector(accu(to_integer(unsigned(din.imm(3 downto 0)))));
	dout.dm_data <= rddata((to_integer(unsigned(din.imm(3 downto 0)))));
	rdaddr <= din.dm_addr;
	-- address for the write needs one cycle delay
	wraddr <= wraddr_dly;
	
	
process(din, rddata)
begin
	if din.dec.sel_imm='1' then
		for i in (stream-1) downto 0 loop
			opd(i) <= unsigned(din.imm);
		end loop;
	else
		-- a MUX for IO will be added
		for i in (stream-1) downto 0 loop
			opd(i) <= unsigned(rddata(i));
		end loop;
	end if;
end process;

-- that's the ALU	
process(din, accu, opd, log, arith, ioin)
begin
	if din.dec.add_sub='0' then
		for i in (stream-1) downto 0 loop
			arith(i) <= accu(i) + opd(i);
		end loop;
	else
		for i in (stream-1) downto 0 loop
			arith(i) <= accu(i) - opd(i);
		end loop;
	end if;

	case din.dec.op is
		when op_ld =>
			for i in (stream-1) downto 0 loop
				log(i) <= opd(i);
			end loop;
		when op_and =>
			for i in (stream-1) downto 0 loop
				log(i) <= accu(i) and opd(i);
			end loop;
		when op_or =>
			for i in (stream-1) downto 0 loop
				log(i) <= accu(i) or opd(i);
			end loop;
		when op_xor =>
			for i in (stream-1) downto 0 loop
				log(i) <= accu(i) xor opd(i);
			end loop;
		when others =>
			null;
	end case;
	
	if din.dec.log_add='0' then
		if din.dec.shr='1' then
			for i in (stream-1) downto 0 loop
				a_mux(i) <= '0' & accu(i)(15 downto 1);
			end loop;
		else
			if din.dec.inp='1' then
				for i in (stream-1) downto 0 loop
					a_mux(i) <= unsigned(ioin.rddata);
				end loop;
			else
				for i in (stream-1) downto 0 loop
					a_mux(i) <= log(i);
				end loop;
			end if;
		end if;
	else
		for i in (stream-1) downto 0 loop	
			a_mux(i) <= arith(i);
		end loop;
	end if;
		
end process;

-- a MUX between 'normal' data and the PC for jal
process(din, accu, pc_dly)
begin
	if din.dec.jal='1' then
		for i in (stream-1) downto 0 loop
			wrdata(i)(IM_BITS-1 downto 0) <= pc_dly;
			wrdata(i)(15 downto IM_BITS) <= (others => '0');
		end loop;
	else
		for i in (stream-1) downto 0 loop
			wrdata(i) <= std_logic_vector(accu(i));
			end loop;
	end if;
end process;	


process(clk, reset)
begin
	if reset='1' then
		accu <= (others => (others => '0'));
--		dout.outp <= (others => '0');
	elsif rising_edge(clk) then
		if din.dec.al_ena = '1' then
			for i in (stream-1) downto 0 loop
				accu(i)(7 downto 0) <= a_mux(i)(7 downto 0);
			end loop;
		end if;
		if din.dec.ah_ena = '1' then
			for i in (stream-1) downto 0 loop
				accu(i)(15 downto 8) <= a_mux(i)(15 downto 8);
			end loop;
		end if;
		wraddr_dly <= din.dm_addr;
		pc_dly <= din.pc;
		-- a simple output port for the hello world example
---             if din.dec.outp='1' then
---                     dout.outp <= std_logic_vector(accu);
---             end if;
	end if;
end process;

-- the data memory (DM)
-- read during write is usually undefined in an FPGA,
-- but that is not modelled
process (clk)
begin
	if rising_edge(clk) then
		-- is store overloaded?
		-- now we have only 'register' read and write
		if din.dec.store='1' then
		for i in (stream-1) downto 0 loop
			dm(i)(to_integer(unsigned(wraddr))) <= wrdata(i);
		end loop;
		end if;
		for i in (stream-1) downto 0 loop
			rddata(i) <= dm(i)(to_integer(unsigned(rdaddr)));
		end loop;
		
	end if;
end process;

	
end rtl;
